module axi4_wrapper #
(
	parameter ;
)(
	input ;
	output ;
);


 endmodule
